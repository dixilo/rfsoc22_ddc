`timescale 1 ps / 1 ps

module system_top(
    input  wire        adc0_clk_clk_n,
    input  wire        adc0_clk_clk_p,
    input  wire        adc2_clk_clk_n,
    input  wire        adc2_clk_clk_p,
    input  wire        dac0_clk_clk_n,
    input  wire        dac0_clk_clk_p,
    input  wire        dac1_clk_clk_n,
    input  wire        dac1_clk_clk_p,
    output wire        ddr4_pl_act_n,
    output wire [16:0] ddr4_pl_adr,
    output wire [1:0]  ddr4_pl_ba,
    output wire [0:0]  ddr4_pl_bg,
    output wire [0:0]  ddr4_pl_ck_c,
    output wire [0:0]  ddr4_pl_ck_t,
    output wire [0:0]  ddr4_pl_cke,
    output wire [0:0]  ddr4_pl_cs_n,
    inout  wire [7:0]  ddr4_pl_dm_n,
    inout  wire [63:0] ddr4_pl_dq,
    inout  wire [7:0]  ddr4_pl_dqs_c,
    inout  wire [7:0]  ddr4_pl_dqs_t,
    output wire [0:0]  ddr4_pl_odt,
    output wire        ddr4_pl_reset_n,
    input  wire        dp_aux_data_in,
    output wire [0:0]  dp_aux_data_oe,
    output wire        dp_aux_data_out,
    input  wire        dp_hot_plug_detect,
    output wire [0:0]  lmk_reset,
    input  wire [0:0]  pl_sysref_n,
    input  wire [0:0]  pl_sysref_p,
    input  wire [0:0]  sys_clk_ddr4_clk_n,
    input  wire [0:0]  sys_clk_ddr4_clk_p,
    input  wire        sysref_in_diff_n,
    input  wire        sysref_in_diff_p,
    input  wire        vin0_01_v_n,
    input  wire        vin0_01_v_p,
    input  wire        vin2_01_v_n,
    input  wire        vin2_01_v_p,
    output wire        vout00_v_n,
    output wire        vout00_v_p,
    output wire        vout10_v_n,
    output wire        vout10_v_p);

    
    wire sysref_int;

    IBUFDS #(
        .DQS_BIAS("FALSE")
    )
    IBUFDS_inst (
        .O(sysref_int),
        .I(pl_sysref_p),
        .IB(pl_sysref_n))
    );

    module system_wrapper(
        .adc0_clk_clk_n(adc0_clk_clk_n),
        .adc0_clk_clk_p(adc0_clk_clk_p),
        .adc2_clk_clk_n(adc2_clk_clk_n),
        .adc2_clk_clk_p(adc2_clk_clk_p),
        .dac0_clk_clk_n(dac0_clk_clk_n),
        .dac0_clk_clk_p(dac0_clk_clk_p),
        .dac1_clk_clk_n(dac1_clk_clk_n),
        .dac1_clk_clk_p(dac1_clk_clk_p),
        .ddr4_pl_act_n(ddr4_pl_act_n),
        .ddr4_pl_adr(ddr4_pl_adr),
        .ddr4_pl_ba(ddr4_pl_ba),
        .ddr4_pl_bg(ddr4_pl_bg),
        .ddr4_pl_ck_c(ddr4_pl_ck_c),
        .ddr4_pl_ck_t(ddr4_pl_ck_t),
        .ddr4_pl_cke(ddr4_pl_cke),
        .ddr4_pl_cs_n(ddr4_pl_cs_n),
        .ddr4_pl_dm_n(ddr4_pl_dm_n),
        .ddr4_pl_dq(ddr4_pl_dq),
        .ddr4_pl_dqs_c(ddr4_pl_dqs_c),
        .ddr4_pl_dqs_t(ddr4_pl_dqs_t),
        .ddr4_pl_odt(ddr4_pl_odt),
        .ddr4_pl_reset_n(ddr4_pl_reset_n),
        .dp_aux_data_in(dp_aux_data_in),
        .dp_aux_data_oe(dp_aux_data_oe),
        .dp_aux_data_out(dp_aux_data_out),
        .dp_hot_plug_detect(dp_hot_plug_detect),
        .lmk_reset(lmk_reset),
        .pl_sysref_in(sysref_int),
        .sys_clk_ddr4_clk_n(sys_clk_ddr4_clk_n),
        .sys_clk_ddr4_clk_p(sys_clk_ddr4_clk_p),
        .sysref_in_diff_n(sysref_in_diff_n),
        .sysref_in_diff_p(sysref_in_diff_p),
        .vin0_01_v_n(vin0_01_v_n),
        .vin0_01_v_p(vin0_01_v_p),
        .vin2_01_v_n(vin2_01_v_n),
        .vin2_01_v_p(vin2_01_v_p),
        .vout00_v_n(vout00_v_n),
        .vout00_v_p(vout00_v_p),
        .vout10_v_n(vout10_v_n),
        .vout10_v_(vout10_v_)
    );
